//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Apr 07 22:42:47 2024
`default_nettype wire
module bootrom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hC20C020029CA10D37848A101DB000DD29108D3004001A83E00D3883E04D39B3E;
defparam prom_inst_0.INIT_RAM_01 = 256'hDCF03100D3063EC9000039C3002EC2BC2370E03EC000210039C3001DC204001D;
defparam prom_inst_0.INIT_RAM_02 = 256'hC4E911062A210272CD76FB0045C20481362C7119712D0491CD6A60FF0E000911;
defparam prom_inst_0.INIT_RAM_03 = 256'h00ACCAEFFE06DBCAFBFEDEF73ADCF432DCF132C33EE500B5210607CD0706083E;
defparam prom_inst_0.INIT_RAM_04 = 256'h02B8CA012FCD04E9C204AACD00A6CAD7FE00A0CACFFE009ACAE7FE0397CAF7FE;
defparam prom_inst_0.INIT_RAM_05 = 256'h72CD76FB00D3033E00F9CD0397C30246C200FECD013AC200D0CD0766C20753CD;
defparam prom_inst_0.INIT_RAM_06 = 256'hE3E307D37904D38B3E4FE0F607DB040600BCC300D33D00CBC2073E08E6790302;
defparam prom_inst_0.INIT_RAM_07 = 256'h823EC904D39B3EB700DBC20500F9CA08E62F05DB07D3A17F3E00F9CA08E605DB;
defparam prom_inst_0.INIT_RAM_08 = 256'h7FE6780125C2AAFE06DB07D3FF3E0125C255FE06DB07D3FE3E05D378FF0604D3;
defparam prom_inst_0.INIT_RAM_09 = 256'h02082105FDCDC9B919DBE3E34F19D30B3EC9B7AF0104FA4720D678012DC3573C;
defparam prom_inst_0.INIT_RAM_0A = 256'h1FE606DB0149C240FE70E605DB0A064F1FE607DB00F9CDDCF522014921DCF222;
defparam prom_inst_0.INIT_RAM_0B = 256'hFE70E605DB0149CA15FA1605D3AF06D37904D3983E4706DB0153C2050149C2B9;
defparam prom_inst_0.INIT_RAM_0C = 256'hC21DDCF4C2AAFE019ECA55FEDCF1CD083E031E0149C2E0E67800F9CD0177C270;
defparam prom_inst_0.INIT_RAM_0D = 256'h01F3CAB77EF50424CD462B57DCF4C2BE2B7EDEF12101A2C2B77E5F0424CD018F;
defparam prom_inst_0.INIT_RAM_0E = 256'h69C101D3C2150C2377AE0A027E207E1123C5D501B7C2BB7E23F14F8787878787;
defparam prom_inst_0.INIT_RAM_0F = 256'hCA03C9CD0000C23C01B7CA93F1C901B7C201FE7A01B7CA03C9CDD1730491CD60;
defparam prom_inst_0.INIT_RAM_10 = 256'hBB0000CA40FEA205DB601EC9D10215CD023DCCFFFE7016D501B7C315041D0000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0215CDC9F100F9CD022DC2BAA205DB0238CA1D05D3AF04D39A3EF506DB0217C2;
defparam prom_inst_0.INIT_RAM_12 = 256'h03230206DB05D37C07D37D4D45800021D10602CDD5873E06A721C9023DC2E6FE;
defparam prom_inst_0.INIT_RAM_13 = 256'h0CD37E02D3780F06E5C5F502A821C90268C2BA7C240386CD0000210255C2BA78;
defparam prom_inst_0.INIT_RAM_14 = 256'hD3AF00D3883EDEF73202DB03D3FD3E00D38A3E027AF20CD3051D0CD3230CD31C;
defparam prom_inst_0.INIT_RAM_15 = 256'h010021000032C33E80802D2D80802D2D80802D2D80802D2DC9F1C1E103D33D02;
defparam prom_inst_0.INIT_RAM_16 = 256'hC20343CDDFE021010E036ACD1BD3AF0376CDDED032343E0600CD069321000122;
defparam prom_inst_0.INIT_RAM_17 = 256'h47DFE43A120000C29602ECC2780D1B23127E4786663E1F0EDEF111DFE0210000;
defparam prom_inst_0.INIT_RAM_18 = 256'h76CDDED03204EEDED03A0305C2B9063E0C0331CA050000C20343CD010E008021;
defparam prom_inst_0.INIT_RAM_19 = 256'hC205240386CD470707DFE43A0100210303C3036ACD1BD3583E0303CA04E67A03;
defparam prom_inst_0.INIT_RAM_1A = 256'h7718DB0356CA92A31BDB0350D20F1BDB1BD3803E01031119D379036ACDC9033A;
defparam prom_inst_0.INIT_RAM_1B = 256'h0377DA7A071BDB1CD357C9036ADA0F1BDB1CD3DED03AC99CE61BDB2B0356F223;
defparam prom_inst_0.INIT_RAM_1C = 256'h3E0602CD0D3E066221C9E1C1038DC20D2C7E36080E0491CDC5E5C000FE7D77C9;
defparam prom_inst_0.INIT_RAM_1D = 256'h03B3DABC03F9CD67825F1FB75703F9CDDCF522039721DCF222044821DEF63211;
defparam prom_inst_0.INIT_RAM_1E = 256'h5F10E601DBD5C9A703CFC281FE23C8A77E0491CD60002E018FC30C1EDEF63282;
defparam prom_inst_0.INIT_RAM_1F = 256'hB74703DACDD5E5C9D187877A03EBCABB1410E601DB01165F03E0CABB10E601DB;
defparam prom_inst_0.INIT_RAM_20 = 256'h290407C21503FBD2B993780417D2905FD1195F0016D503DACD20160000214F1F;
defparam prom_inst_0.INIT_RAM_21 = 256'h9696782B042FC20D083E47802377DCF1CDFF3E002301E5DED021D5C5C9E1D17C;
defparam prom_inst_0.INIT_RAM_22 = 256'h1779070707070452CABB10E601DB5F10E601DB57000ED5C5C9C1D10429C2E17E;
defparam prom_inst_0.INIT_RAM_23 = 256'h3E044DC219FE0484C3DEF432AF047AC2E6FE790486F2B77A0464C23DDEF63A4F;
defparam prom_inst_0.INIT_RAM_24 = 256'hC685821F5770E61F7C6F0707077DD5C9C1D1A9DEF43A044DC2150916DEF432FF;
defparam prom_inst_0.INIT_RAM_25 = 256'h003E0553CDDED4323CDED332DED232AFDED522FF0021C9D167C0C61FE67C6F18;
defparam prom_inst_0.INIT_RAM_26 = 256'h534F00C9B7E13D04CCC20D231304DAC2003EBE1A0C0E04DD11E5FF002104DBC2;
defparam prom_inst_0.INIT_RAM_27 = 256'hCAB77E100EFF102144DED5220100210602CD8C3E067C214D4F43202020202020;
defparam prom_inst_0.INIT_RAM_28 = 256'hC3190010110522CA04C6CD04FDC20D230000C2B7DED23A4704C6780529CD0522;
defparam prom_inst_0.INIT_RAM_29 = 256'hF1DED232FF3E053FCA0553CDF5DED432013EDED332E5F50268C30100215004FB;
defparam prom_inst_0.INIT_RAM_2A = 256'hF3058CCDDED02239000021D5C5C9F1E10530C209FE3CDED52219008011DED52A;
defparam prom_inst_0.INIT_RAM_2B = 256'h10D3003E4F0569C20D237223738283D1237223738283D1200EAFDED52AF910D3;
defparam prom_inst_0.INIT_RAM_2C = 256'hFE2FDED33AEB0595C23D19040021FF8011DED43AC9C1D105D7CD79FBF9DED02A;
defparam prom_inst_0.INIT_RAM_2D = 256'h3AC9C1B1103E4FC50CE60707070719002E7D67FCE607076F04D610D605A6D2FC;
defparam prom_inst_0.INIT_RAM_2E = 256'hDED02239000021D5F5C91C3E6F85873DDED43A6784F03E2929292900266FDED3;
defparam prom_inst_0.INIT_RAM_2F = 256'h06B521C9FF3EC89505FAC2BCF1D1EBFBF9DED02A10D3003ED1F910D3F305BFCD;
defparam prom_inst_0.INIT_RAM_30 = 256'h0D2313127E061EF2B7DCF73A13127ED54F7FE6DCF73ADCF732D8E21102068A3E;
defparam prom_inst_0.INIT_RAM_31 = 256'h181818181818DB1B1A9C1A1B1BDBF3DBDBF3DBDBDBF3C9060AC20514D10611C2;
defparam prom_inst_0.INIT_RAM_32 = 256'h1696D6D6DF83E3B6B6B7B6B6B6E3C061616D6DC1010073DBDBDBDBDBDB737E5A;
defparam prom_inst_0.INIT_RAM_33 = 256'h9280FF0FFE0301FFFF3723F7FF03FDD5FC7FC080FFFFECC4EFFFC0BFAB3F96D6;
defparam prom_inst_0.INIT_RAM_34 = 256'h7F7FFFFF8181FFFCFCFFFEFEFF014901490149014901FFF0FF80928092809280;
defparam prom_inst_0.INIT_RAM_35 = 256'h83C1200704E407010F20C154FF03C603FF5455FFC0C7C0FF55FFFFFEFF3F3FFF;
defparam prom_inst_0.INIT_RAM_36 = 256'h823E05FDCD80FF80FF80FF80FF8001FF01FF01FF01FF018304E02027E080F004;
defparam prom_inst_0.INIT_RAM_37 = 256'hCD63071CCD0000C2AAFE7B071CCD0000C255FE7B071CCD4F6FAF05D3103E04D3;
defparam prom_inst_0.INIT_RAM_38 = 256'h06DB0016C7C8B97B071CCD0705C2B87C230382CD4FAB7973071CCD47837C071C;
defparam prom_inst_0.INIT_RAM_39 = 256'hAF00165FB3070707070FE606DB073FC3145F0FE606DB0733C2A77A071ECA20E6;
defparam prom_inst_0.INIT_RAM_3A = 256'hFEC0E657DBC8050F065FD3803EC9071EC2A77A05D3103E0742C220E606DB05D3;
defparam prom_inst_0.INIT_RAM_3B = 256'h043A07D5CD0000CAE5FEE4043A0792CD013E0602CD893E06C921C9B70759C240;
defparam prom_inst_0.INIT_RAM_3C = 256'h53D37D2C002E0026E000114F873CC90268CD57848787E4043AE4002A0792CDE4;
defparam prom_inst_0.INIT_RAM_3D = 256'hCD58DB07EFCD50DB0006E107D7CD5826E557D3203E52D33C55D354D3AF56D37C;
defparam prom_inst_0.INIT_RAM_3E = 256'hCABCD9E657DB2006C55026079AC324079CC2BDE0803A07D5CA0D07B8C20507EF;
defparam prom_inst_0.INIT_RAM_3F = 256'hC9E1EBE4002AE5C080FE7BC0E4FE7A1312C9C1C707DAC2B1780B07DAC22D07ED;

endmodule //bootrom
